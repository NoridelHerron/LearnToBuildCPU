`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Create Date: 08/16/2025 07:38:43 AM
// Module Name: rom
// Created by: Noridel Herron
//////////////////////////////////////////////////////////////////////////////////
`include "constant_def.vh"

module rom_v ( 
       input  wire        clk,
       input  wire [9:0]  addr,    // PC >> 2 for word indexing
       output reg  [31:0] instr
    );
    reg [31:0] rom [0:1023];
    reg [14:0] temp_reg;
    /*
    function [14:0] generate_registers;
        input integer type_sel;
        input reg [4:0] rd;
        reg [14:0] rand_reg;
        
         begin
            case (type_sel) // rd = rand_reg[14:10], rs2= rand_reg[9:5], rs1 = rand_reg[4:0]
               // Case 0-2 will help generate hazard later
               0 : begin 
                    rand_reg[14:10] = $urandom_range(0, 31); 
                    rand_reg[9:5]   = rd; 
                    rand_reg[4:0]   = $urandom_range(0, 31);
               end 
               
               1 : begin 
                    rand_reg[14:10] = $urandom_range(0, 31); 
                    rand_reg[9:5]   =  $urandom_range(0, 31); 
                    rand_reg[4:0]   = rd; 
               end 
               
               2 : begin 
                    rand_reg[14:10] = $urandom_range(0, 31); 
                    rand_reg[9:5]   = rd; 
                    rand_reg[4:0]   = rd; 
               end 
               
               3 : begin 
                    rand_reg[14:10] = $urandom_range(0, 31); 
                    rand_reg[9:5]   =  $urandom_range(0, 31); 
                    rand_reg[4:0]   = $urandom_range(0, 31); 
               end 
               
               default : begin 
                    rand_reg[14:10] = $urandom_range(1, 31); 
                    rand_reg[9:5]   =  $urandom_range(1, 31); 
                    rand_reg[4:0]   = $urandom_range(1, 31); 
               end 
            endcase
        generate_registers = rand_reg;
        end
    endfunction
    
    function [31:0] generate_instruction;
        input integer type_sel;
        input [14:0] registers;
        reg [2:0]  funct3;
        reg [6:0]  funct7;
        reg [11:0] imm12;  // 12-bit immediate // divisible by 4
        reg [19:0] imm20;  // 20-bit immediate // divisible by 4
        reg [31:0] instr;

        begin
            funct3 = $urandom_range(0, 7);
            funct7 = $urandom_range(0, 127);

            case (type_sel)
            
                //==== R-type logic (e.g., add, sub, srl, sra) ====
                0: begin
                    if (funct3 == `F3_ADD_SUB || funct3 == `F3_SRL_SRA) begin
                        funct7 = $urandom_range(0, 1) ? 7'd0 : 7'd32;  // ADD/SRL or SUB/SRA
                    end else begin
                        funct7 = 7'd0; // other R-type
                    end
                    instr = {funct7, registers[9:5], registers[4:0], funct3, registers[14:0], `R_TYPE};
                end

                //==== I-type Immediate ====
                1: begin
                    imm12 = {funct7, registers[9:5]} * 4; 
                    instr = {imm12, registers[4:0], funct3, registers[14:0], `I_IMM};
                end

                // ==== Load (e.g., LW) ====
                2: begin
                    funct3 = `F3_LW; // Force LW
                    imm12 = {funct7, registers[9:5]} * 4; 
                    instr = {imm12, registers[4:0], funct3, registers[14:0], `I_LOAD};
                end
                
                // ===== S-type logic (e.g., store) ===
                3: begin
                    funct3 = `F3_SW; // Force LW
                    imm12 = {funct7, registers[9:5]} * 4; 
                    instr = {imm12[11:5], registers[9:5], registers[4:0], funct3, imm12[4:0], `S_TYPE};
                end
                
                //==== B-type logic (e.g., beq) ====
                4: begin
                    case (funct3)
                        0: funct3 = `BEQ;
                        1: funct3 = `BNE;
                        4: funct3 = `BLT;
                        5: funct3 = `BGE;
                        6: funct3 = `BLTU;
                        7: funct3 = `BGEU;
                        default: funct3 = $urandom_range(4, 7);
                    endcase
                    imm12 = {funct7, registers[9:5]} * 4; 
                    instr = {imm12[11], imm12[9:4], registers[9:5], registers[4:0], 
                             funct3, imm12[3:0], imm12[10], `B_TYPE};
                end

                // ==== JAL Logic ====
                5: begin
                    imm20 = {funct7, registers[9:5], registers[4:0], funct3}; // 20-bit signed immediate
                    instr = {
                                imm20[19],       // bit 31
                                imm20[9:0],      // bits 30:21
                                imm20[10],       // bit 20
                                imm20[18:11],    // bits 19:12
                                registers[14:0], // bits 11:7
                                `J_JAL     // bits 6:0
                            };
                end

                //==== Default (NOP) ====
                default: instr = 32'h00000013;

            endcase

            generate_instruction = instr;
        end
    endfunction
    
    integer i;
    
    initial begin
        $display("ROM STARTED");
        for (i = 0; i < 1024; i = i + 1) begin
            temp_reg = generate_registers ($urandom_range(3, 5), 5'b0);
            rom[i] = generate_instruction($urandom_range(0, 5), temp_reg);
            $display("ROM[%0d] = %h", i, rom[i]);
        end 
    end
    */
    initial begin
        rom[0] = 32'h008C2503;
rom[1] = 32'h6A0930EF;
rom[2] = 32'hBBCCA223;
rom[3] = 32'h5A131CE3;
rom[4] = 32'hF0491C6F;
rom[5] = 32'h080C4863;
rom[6] = 32'h01721FB3;
rom[7] = 32'h6A3A5463;
rom[8] = 32'h14C5A823;
rom[9] = 32'h01CD6733;
rom[10] = 32'h004213B3;
rom[11] = 32'h532BEE6F;
rom[12] = 32'h0011C9B3;
rom[13] = 32'h03342E23;
rom[14] = 32'hA60F2E23;
rom[15] = 32'h6ED68CE3;
rom[16] = 32'h68302023;
rom[17] = 32'h17096F93;
rom[18] = 32'h052900EF;
rom[19] = 32'h2571AC23;
rom[20] = 32'h695B7C63;
rom[21] = 32'h01E5CA33;
rom[22] = 32'hDFBBAA23;
rom[23] = 32'h4B57A223;
rom[24] = 32'h7B83EB13;
rom[25] = 32'h0002A503;
rom[26] = 32'h002A8EB3;
rom[27] = 32'h00AAE5B3;
rom[28] = 32'h6D09916F;
rom[29] = 32'h55972A23;
rom[30] = 32'h0181A003;
rom[31] = 32'hDDAA2823;
rom[32] = 32'h0104FBB3;
rom[33] = 32'hE2411393;
rom[34] = 32'h0105A983;
rom[35] = 32'h7F3D7863;
rom[36] = 32'hC824AC23;
rom[37] = 32'h83F64B6F;
rom[38] = 32'h46EAA823;
rom[39] = 32'h48D984E3;
rom[40] = 32'hF5F6A423;
rom[41] = 32'h0060E9B3;
rom[42] = 32'h01442783;
rom[43] = 32'h063F9063;
rom[44] = 32'h104A2B93;
rom[45] = 32'h011163B3;
rom[46] = 32'h01082883;
rom[47] = 32'h44656C63;
rom[48] = 32'hCD08AD93;
rom[49] = 32'h00C62A03;
rom[50] = 32'h000AA203;
rom[51] = 32'h5DB14CE3;
rom[52] = 32'h23DBA623;
rom[53] = 32'h114CAA23;
rom[54] = 32'h00812303;
rom[55] = 32'h0043E133;
rom[56] = 32'hFE91A023;
rom[57] = 32'h31BD08E3;
rom[58] = 32'h1054626F;
rom[59] = 32'h01CD2983;
rom[60] = 32'h008AA803;
rom[61] = 32'hBCA8916F;
rom[62] = 32'h0049A483;
rom[63] = 32'h1A322E23;
rom[64] = 32'h36E9C4E3;
rom[65] = 32'h004A6FB3;
rom[66] = 32'h018DAA03;
rom[67] = 32'h92CEB893;
rom[68] = 32'h7D097713;
rom[69] = 32'h7D91D8E3;
rom[70] = 32'h09081893;
rom[71] = 32'h00CC2B83;
rom[72] = 32'h01931633;
rom[73] = 32'h008AAA03;
rom[74] = 32'h31089513;
rom[75] = 32'h47549863;
rom[76] = 32'hF695A223;
rom[77] = 32'h8F079093;
rom[78] = 32'h01A2F1B3;
rom[79] = 32'h014D2D03;
rom[80] = 32'h0E13CEEF;
rom[81] = 32'h00C8AC03;
rom[82] = 32'h01FF20B3;
rom[83] = 32'h052CA06F;
rom[84] = 32'h00B6E9B3;
rom[85] = 32'h7BE404E3;
rom[86] = 32'h019592B3;
rom[87] = 32'h41895913;
rom[88] = 32'h9D8E83EF;
rom[89] = 32'h00092E03;
rom[90] = 32'h783F2423;
rom[91] = 32'h01052103;
rom[92] = 32'hD712A623;
rom[93] = 32'hC582C1EF;
rom[94] = 32'h4669DCE3;
rom[95] = 32'hF8D710EF;
rom[96] = 32'h01C7AE83;
rom[97] = 32'h46A4E463;
rom[98] = 32'hC3453193;
rom[99] = 32'h01CCAB83;
rom[100] = 32'hB88E2423;
rom[101] = 32'h00F1AB33;
rom[102] = 32'h40895F93;
rom[103] = 32'hC2BE616F;
rom[104] = 32'hCDA0A223;
rom[105] = 32'h4B0E1463;
rom[106] = 32'h00A7F4B3;
rom[107] = 32'h2D3110E3;
rom[108] = 32'h014CA703;
rom[109] = 32'h888AE093;
rom[110] = 32'h01BA4433;
rom[111] = 32'h01CEA583;
rom[112] = 32'h4709E66F;
rom[113] = 32'h01492403;
rom[114] = 32'h004B01B3;
rom[115] = 32'h00F282EF;
rom[116] = 32'h8ACB8DEF;
rom[117] = 32'h6C9A9463;
rom[118] = 32'h4319A623;
rom[119] = 32'h2AB42223;
rom[120] = 32'h010CA783;
rom[121] = 32'h20638CE3;
rom[122] = 32'h010DA483;
rom[123] = 32'h010BAB83;
rom[124] = 32'h69D00CE3;
rom[125] = 32'h002608B3;
rom[126] = 32'h01524AB3;
rom[127] = 32'h00DFF733;
rom[128] = 32'h00CDAD83;
rom[129] = 32'h2BFFA023;
rom[130] = 32'hA2F20EEF;
rom[131] = 32'h6EDD6B6F;
rom[132] = 32'h49659463;
rom[133] = 32'h017723B3;
rom[134] = 32'h0106D913;
rom[135] = 32'h080D8693;
rom[136] = 32'h00FB2C33;
rom[137] = 32'h2C0F0113;
rom[138] = 32'h18887CE3;
rom[139] = 32'h177D5C63;
rom[140] = 32'h18925863;
rom[141] = 32'h5093C2EF;
rom[142] = 32'h01A4A9B3;
rom[143] = 32'hE5CCC9EF;
rom[144] = 32'h45AA2823;
rom[145] = 32'h61C5CA13;
rom[146] = 32'h01C82C03;
rom[147] = 32'hDC94236F;
rom[148] = 32'h63B584E3;
rom[149] = 32'h01A7E1B3;
rom[150] = 32'hC4D82623;
rom[151] = 32'h00837C13;
rom[152] = 32'hC02B87EF;
rom[153] = 32'hD8899C13;
rom[154] = 32'hA0862A6F;
rom[155] = 32'h0BBE2823;
rom[156] = 32'h7C4C9613;
rom[157] = 32'h6A6804E3;
rom[158] = 32'h00C9AC03;
rom[159] = 32'h8C069E93;
rom[160] = 32'hA69109EF;
rom[161] = 32'hD5DDA823;
rom[162] = 32'h39ED876F;
rom[163] = 32'h3769EC63;
rom[164] = 32'h59920463;
rom[165] = 32'h3BB71B6F;
rom[166] = 32'h01605633;
rom[167] = 32'h9AB7A023;
rom[168] = 32'h40805493;
rom[169] = 32'h486179EF;
rom[170] = 32'h7B0CBE13;
rom[171] = 32'hB476426F;
rom[172] = 32'h8BCFC893;
rom[173] = 32'h34E22A23;
rom[174] = 32'h0124FE33;
rom[175] = 32'h014A4133;
rom[176] = 32'h003E1063;
rom[177] = 32'h00CC45B3;
rom[178] = 32'hC757A623;
rom[179] = 32'h443FF0E3;
rom[180] = 32'hC9612823;
rom[181] = 32'hF71C2623;
rom[182] = 32'h05EF2223;
rom[183] = 32'h0184A503;
rom[184] = 32'h4E19AFEF;
rom[185] = 32'h004CA903;
rom[186] = 32'hFB2BA26F;
rom[187] = 32'h0082A883;
rom[188] = 32'h61E784E3;
rom[189] = 32'h643C5CE3;
rom[190] = 32'h41288333;
rom[191] = 32'hE1BA2623;
rom[192] = 32'h0110BB33;
rom[193] = 32'h014DA9B3;
rom[194] = 32'h95E1A623;
rom[195] = 32'h40BB5B33;
rom[196] = 32'h8C0C9F13;
rom[197] = 32'h01462E83;
rom[198] = 32'h01D71CB3;
rom[199] = 32'hBC32A223;
rom[200] = 32'h41085393;
rom[201] = 32'h0081AA03;
rom[202] = 32'h000DAE03;
rom[203] = 32'h09539CE3;
rom[204] = 32'h52026893;
rom[205] = 32'h8517A023;
rom[206] = 32'h0046BBB3;
rom[207] = 32'h008F2B03;
rom[208] = 32'hBA811C13;
rom[209] = 32'h98B52623;
rom[210] = 32'h01C92783;
rom[211] = 32'h6A84DE6F;
rom[212] = 32'h62FD7863;
rom[213] = 32'h738B7293;
rom[214] = 32'h024F8C63;
rom[215] = 32'hFCB72623;
rom[216] = 32'h01452EB3;
rom[217] = 32'h8043CC13;
rom[218] = 32'h0045AE03;
rom[219] = 32'h64402413;
rom[220] = 32'h3B8963EF;
rom[221] = 32'h5FFC846F;
rom[222] = 32'h018E45B3;
rom[223] = 32'hA08B8F93;
rom[224] = 32'hF436C5EF;
rom[225] = 32'h01CE13B3;
rom[226] = 32'h34019193;
rom[227] = 32'h9758A223;
rom[228] = 32'h0188F933;
rom[229] = 32'h298317EF;
rom[230] = 32'h0041AE83;
rom[231] = 32'h67BDD26F;
rom[232] = 32'h01C02E83;
rom[233] = 32'h3019816F;
rom[234] = 32'h65C564E3;
rom[235] = 32'hA5E0AE23;
rom[236] = 32'hA94D2A23;
rom[237] = 32'h01852C83;
rom[238] = 32'h110BAC23;
rom[239] = 32'h32AC1063;
rom[240] = 32'hF8CF3F13;
rom[241] = 32'h00CD5513;
rom[242] = 32'h71567CE3;
rom[243] = 32'h400D5733;
rom[244] = 32'hE4FEF6EF;
rom[245] = 32'h00472983;
rom[246] = 32'hBC30A023;
rom[247] = 32'h0132B4B3;
rom[248] = 32'h6F141C63;
rom[249] = 32'hA8F0CCEF;
rom[250] = 32'hA785F593;
rom[251] = 32'h364C6893;
rom[252] = 32'h00CCAB03;
rom[253] = 32'h00C69C33;
rom[254] = 32'h45ECC863;
rom[255] = 32'h2B4FE863;
rom[256] = 32'h08046A93;
rom[257] = 32'h018CB6B3;
rom[258] = 32'h3BFFE0E3;
rom[259] = 32'h0DB5A023;
rom[260] = 32'h5881B393;
rom[261] = 32'h3E21F4EF;
rom[262] = 32'h2552D863;
rom[263] = 32'h00CB2683;
rom[264] = 32'h1C64B06F;
rom[265] = 32'h01432603;
rom[266] = 32'h4018D5B3;
rom[267] = 32'h009AECB3;
rom[268] = 32'h24419793;
rom[269] = 32'h01092B83;
rom[270] = 32'h77E74863;
rom[271] = 32'h00082E03;
rom[272] = 32'h7E1AAC23;
rom[273] = 32'h39D3A823;
rom[274] = 32'h01831033;
rom[275] = 32'h651248E3;
rom[276] = 32'hC81A2823;
rom[277] = 32'hF54A6F13;
rom[278] = 32'h1FECADEF;
rom[279] = 32'hADF9B26F;
rom[280] = 32'hA378EC6F;
rom[281] = 32'h03E000E3;
rom[282] = 32'h4816D4E3;
rom[283] = 32'h018BA983;
rom[284] = 32'h49BCD063;
rom[285] = 32'hF0443413;
rom[286] = 32'h07ADCEEF;
rom[287] = 32'hED922023;
rom[288] = 32'h113EAE23;
rom[289] = 32'h00092503;
rom[290] = 32'hD689A023;
rom[291] = 32'h6E5004E3;
rom[292] = 32'h00062F83;
rom[293] = 32'h49052493;
rom[294] = 32'h01C5A683;
rom[295] = 32'h0007A483;
rom[296] = 32'h843C2223;
rom[297] = 32'h008E2483;
rom[298] = 32'h2E971063;
rom[299] = 32'h00CCF9B3;
rom[300] = 32'h01E19D33;
rom[301] = 32'hF1008393;
rom[302] = 32'h96C3A223;
rom[303] = 32'h01294433;
rom[304] = 32'hDD23D0EF;
rom[305] = 32'hA637E3EF;
rom[306] = 32'h01C0A703;
rom[307] = 32'h00002803;
rom[308] = 32'h00CCBBB3;
rom[309] = 32'h0045FE33;
rom[310] = 32'h3CD80463;
rom[311] = 32'h5C94EC63;
rom[312] = 32'h00DB7BB3;
rom[313] = 32'hB26A14EF;
rom[314] = 32'h54024393;
rom[315] = 32'hED443993;
rom[316] = 32'h6CD50863;
rom[317] = 32'h71802223;
rom[318] = 32'hB17C2023;
rom[319] = 32'h07BCA823;
rom[320] = 32'h01362FB3;
rom[321] = 32'h60AAD463;
rom[322] = 32'h000C2103;
rom[323] = 32'h00CC2903;
rom[324] = 32'h05D58463;
rom[325] = 32'h67889D13;
rom[326] = 32'h561E05EF;
rom[327] = 32'h0112C533;
rom[328] = 32'hC5D6BCEF;
rom[329] = 32'h563FA823;
rom[330] = 32'h4E97D8E3;
rom[331] = 32'hA1C52823;
rom[332] = 32'h2CCBF393;
rom[333] = 32'hAF422613;
rom[334] = 32'h5FB49863;
rom[335] = 32'h010F2903;
rom[336] = 32'h823BB8EF;
rom[337] = 32'h00345F33;
rom[338] = 32'h737C2A23;
rom[339] = 32'h2CC53093;
rom[340] = 32'h018DA703;
rom[341] = 32'h3EA69CE3;
rom[342] = 32'h5C5D2223;
rom[343] = 32'h36F944EF;
rom[344] = 32'h01B5F333;
rom[345] = 32'h0703A223;
rom[346] = 32'h000ADF13;
rom[347] = 32'h001D66B3;
rom[348] = 32'h394E7E13;
rom[349] = 32'h00CCA683;
rom[350] = 32'h65154463;
rom[351] = 32'h470A26EF;
rom[352] = 32'h0C82FA93;
rom[353] = 32'hE444AA23;
rom[354] = 32'hD0AA2C23;
rom[355] = 32'h71CCF193;
rom[356] = 32'h450D9C63;
rom[357] = 32'h52F804E3;
rom[358] = 32'hCA02A823;
rom[359] = 32'h54C89AEF;
rom[360] = 32'h43E52623;
rom[361] = 32'h2BC96463;
rom[362] = 32'h01FB3CB3;
rom[363] = 32'h4101D793;
rom[364] = 32'h24B07463;
rom[365] = 32'h724D246F;
rom[366] = 32'h7B0800E3;
rom[367] = 32'h00CCAA83;
rom[368] = 32'h468668E3;
rom[369] = 32'h101B246F;
rom[370] = 32'h88EEA96F;
rom[371] = 32'h124A3893;
rom[372] = 32'h2E78A423;
rom[373] = 32'hA720A223;
rom[374] = 32'h11A0D8E3;
rom[375] = 32'h0086A783;
rom[376] = 32'h7603E293;
rom[377] = 32'h1079A823;
rom[378] = 32'h6F962E23;
rom[379] = 32'h5C597463;
rom[380] = 32'h00C748B3;
rom[381] = 32'h3B841C93;
rom[382] = 32'h27BC016F;
rom[383] = 32'h01A39933;
rom[384] = 32'h71453313;
rom[385] = 32'hF62E2E23;
rom[386] = 32'h6C0CD86F;
rom[387] = 32'h47E6A023;
rom[388] = 32'h7F3208E3;
rom[389] = 32'h777AFCE3;
rom[390] = 32'h00777333;
rom[391] = 32'h746CA023;
rom[392] = 32'hBF096893;
rom[393] = 32'h418A5A33;
rom[394] = 32'h0149AA83;
rom[395] = 32'h003234B3;
rom[396] = 32'h00191933;
rom[397] = 32'h0EA03D6F;
rom[398] = 32'h007CCC33;
rom[399] = 32'h95642023;
rom[400] = 32'h01032103;
rom[401] = 32'h467EAE23;
rom[402] = 32'h2288A893;
rom[403] = 32'hE644F613;
rom[404] = 32'hB0302C23;
rom[405] = 32'h00CE2583;
rom[406] = 32'h014FA903;
rom[407] = 32'h019E07B3;
rom[408] = 32'h0B4FDC63;
rom[409] = 32'h60CD3E13;
rom[410] = 32'h2DF5976F;
rom[411] = 32'hBE83206F;
rom[412] = 32'hF1044A93;
rom[413] = 32'h5C491E93;
rom[414] = 32'h6B4E8C63;
rom[415] = 32'hAD813D13;
rom[416] = 32'h008B3433;
rom[417] = 32'h00802603;
rom[418] = 32'hE0C0FA93;
rom[419] = 32'h8E955C6F;
rom[420] = 32'h0006AD83;
rom[421] = 32'hECB1A223;
rom[422] = 32'h685BF9EF;
rom[423] = 32'h380FD063;
rom[424] = 32'hB6432393;
rom[425] = 32'h1CA12423;
rom[426] = 32'h71C5FB93;
rom[427] = 32'h014C2503;
rom[428] = 32'h010E27B3;
rom[429] = 32'h01882803;
rom[430] = 32'h80112023;
rom[431] = 32'hD8018313;
rom[432] = 32'h9B8B2623;
rom[433] = 32'h00E18133;
rom[434] = 32'h81098E13;
rom[435] = 32'h43050C93;
rom[436] = 32'h00C22003;
rom[437] = 32'h01F22733;
rom[438] = 32'h008EAC03;
rom[439] = 32'h5A873B6F;
rom[440] = 32'hFEFDA823;
rom[441] = 32'h00032403;
rom[442] = 32'h0164F8B3;
rom[443] = 32'h530AC063;
rom[444] = 32'h0132EA33;
rom[445] = 32'h40B4D4B3;
rom[446] = 32'hE8B6AC6F;
rom[447] = 32'h01C5A283;
rom[448] = 32'h003764B3;
rom[449] = 32'h4C6314E3;
rom[450] = 32'h4A9254E3;
rom[451] = 32'h492514E3;
rom[452] = 32'h41FC86B3;
rom[453] = 32'h0001AA83;
rom[454] = 32'h339557EF;
rom[455] = 32'h01482883;
rom[456] = 32'h66B12C23;
rom[457] = 32'h9597EEEF;
rom[458] = 32'hCD2C2A23;
rom[459] = 32'h41555433;
rom[460] = 32'h0C971E6F;
rom[461] = 32'h67F0D863;
rom[462] = 32'h9032A823;
rom[463] = 32'h001A7E33;
rom[464] = 32'h0050BCB3;
rom[465] = 32'h65700CE3;
rom[466] = 32'h00C26F33;
rom[467] = 32'h12099C63;
rom[468] = 32'h70879CE3;
rom[469] = 32'hDFEA20EF;
rom[470] = 32'h4A962C23;
rom[471] = 32'h770E9D93;
rom[472] = 32'hAE1D2223;
rom[473] = 32'h01C5A083;
rom[474] = 32'h01082403;
rom[475] = 32'h2DC02A23;
rom[476] = 32'h0140F493;
rom[477] = 32'h5FE51AEF;
rom[478] = 32'h0145A603;
rom[479] = 32'hD1282023;
rom[480] = 32'h01C82D83;
rom[481] = 32'h78639063;
rom[482] = 32'h70018593;
rom[483] = 32'h16DF80E3;
rom[484] = 32'hF538186F;
rom[485] = 32'h01F888E3;
rom[486] = 32'h10D1146F;
rom[487] = 32'h011E21B3;
rom[488] = 32'h018308B3;
rom[489] = 32'h0135CDB3;
rom[490] = 32'h9626A223;
rom[491] = 32'h412E00B3;
rom[492] = 32'h00BEBAB3;
rom[493] = 32'h00AA4433;
rom[494] = 32'h65661863;
rom[495] = 32'hB8CF2023;
rom[496] = 32'h654C8713;
rom[497] = 32'h004FDC13;
rom[498] = 32'h57448E93;
rom[499] = 32'h521DCC6F;
rom[500] = 32'h00A5AA33;
rom[501] = 32'hD18EB513;
rom[502] = 32'h00E10CB3;
rom[503] = 32'h37313AEF;
rom[504] = 32'h004DD913;
rom[505] = 32'h2D9BA7EF;
rom[506] = 32'h54E918E3;
rom[507] = 32'h3EB5A823;
rom[508] = 32'h26E5B16F;
rom[509] = 32'h01CE2603;
rom[510] = 32'h6F5139EF;
rom[511] = 32'h00432F33;
rom[512] = 32'h00E868E3;
rom[513] = 32'hBC468E13;
rom[514] = 32'hEB51486F;
rom[515] = 32'h00052E03;
rom[516] = 32'hCE8E1B93;
rom[517] = 32'h3421C36F;
rom[518] = 32'h4A2A98EF;
rom[519] = 32'h6C5EEEEF;
rom[520] = 32'h010C2803;
rom[521] = 32'h00B756B3;
rom[522] = 32'h744E4CE3;
rom[523] = 32'h786B5CE3;
rom[524] = 32'h9F082A93;
rom[525] = 32'h77460013;
rom[526] = 32'h3DB52223;
rom[527] = 32'hE5C9A313;
rom[528] = 32'h225098E3;
rom[529] = 32'h1C3FA423;
rom[530] = 32'hD315A823;
rom[531] = 32'h01C4A483;
rom[532] = 32'hD2523E6F;
rom[533] = 32'h1EB2FC63;
rom[534] = 32'h03C4E26F;
rom[535] = 32'hD7C71713;
rom[536] = 32'h00889633;
rom[537] = 32'h01012883;
rom[538] = 32'hBE232C23;
rom[539] = 32'h1ED423EF;
rom[540] = 32'h3084AE13;
rom[541] = 32'h000FAC03;
rom[542] = 32'h10449CE3;
rom[543] = 32'h21A694E3;
rom[544] = 32'h000D2B03;
rom[545] = 32'h28EBFCE3;
rom[546] = 32'h571F14E3;
rom[547] = 32'h9280AE93;
rom[548] = 32'h466D2C6F;
rom[549] = 32'h42D994E3;
rom[550] = 32'hE34F9913;
rom[551] = 32'hB3932623;
rom[552] = 32'h1E7D8D6F;
rom[553] = 32'h01CD2903;
rom[554] = 32'h00457333;
rom[555] = 32'h01445C6F;
rom[556] = 32'h74C2A423;
rom[557] = 32'h010FA183;
rom[558] = 32'h01CBA783;
rom[559] = 32'h4090AA23;
rom[560] = 32'h255FFDEF;
rom[561] = 32'h0C7BA023;
rom[562] = 32'h122CA023;
rom[563] = 32'h2016DA6F;
rom[564] = 32'h010E2A83;
rom[565] = 32'h00DCF733;
rom[566] = 32'h6AB92423;
rom[567] = 32'h2491DC63;
rom[568] = 32'h74861CE3;
rom[569] = 32'h7EA12C23;
rom[570] = 32'h01CEA333;
rom[571] = 32'h3C3058E3;
rom[572] = 32'h00806033;
rom[573] = 32'h2F61A023;
rom[574] = 32'h00802103;
rom[575] = 32'h657A11EF;
rom[576] = 32'h411F0733;
rom[577] = 32'h15C72E23;
rom[578] = 32'h6ECB8463;
rom[579] = 32'h9C1AA823;
rom[580] = 32'h00472703;
rom[581] = 32'h4DF91463;
rom[582] = 32'h008DA483;
rom[583] = 32'hA600F993;
rom[584] = 32'h0949E493;
rom[585] = 32'h002CD3B3;
rom[586] = 32'h0048A383;
rom[587] = 32'h00C52D03;
rom[588] = 32'h36F694E3;
rom[589] = 32'h0E2B2423;
rom[590] = 32'h53AFAE23;
rom[591] = 32'h01F2AE33;
rom[592] = 32'h0041A883;
rom[593] = 32'h4E416813;
rom[594] = 32'h00822283;
rom[595] = 32'hD35DE26F;
rom[596] = 32'h400F0433;
rom[597] = 32'hA1CB1E93;
rom[598] = 32'h423FE76F;
rom[599] = 32'h000A2883;
rom[600] = 32'h71CED4E3;
rom[601] = 32'hF74FE293;
rom[602] = 32'h00CA2303;
rom[603] = 32'h01062483;
rom[604] = 32'h01062C83;
rom[605] = 32'h05E47063;
rom[606] = 32'hC7CAA223;
rom[607] = 32'h05319DEF;
rom[608] = 32'h5CB68063;
rom[609] = 32'h01881433;
rom[610] = 32'h9DF1F8EF;
rom[611] = 32'h7A834C93;
rom[612] = 32'h5DAAB86F;
rom[613] = 32'h6C7C6BEF;
rom[614] = 32'h958C3B93;
rom[615] = 32'h01271E33;
rom[616] = 32'h3BFA5463;
rom[617] = 32'h0100D113;
rom[618] = 32'h46469E13;
rom[619] = 32'h00C82903;
rom[620] = 32'h4F75AA23;
rom[621] = 32'h515EA823;
rom[622] = 32'h0108AD03;
rom[623] = 32'h01492883;
rom[624] = 32'h0D2A106F;
rom[625] = 32'h0049A803;
rom[626] = 32'h05ABF063;
rom[627] = 32'h1D4A4FEF;
rom[628] = 32'h68FAA623;
rom[629] = 32'h62BAE863;
rom[630] = 32'h000D5C93;
rom[631] = 32'hF3872623;
rom[632] = 32'h2C0074E3;
rom[633] = 32'h413F85B3;
rom[634] = 32'h00B74433;
rom[635] = 32'h40DF8AB3;
rom[636] = 32'h273678E3;
rom[637] = 32'h3F318863;
rom[638] = 32'h46B29463;
rom[639] = 32'h0033A733;
rom[640] = 32'h00911CB3;
rom[641] = 32'h01A27E33;
rom[642] = 32'hF81D7A6F;
rom[643] = 32'h847B446F;
rom[644] = 32'h40CFD7B3;
rom[645] = 32'hB88FAC23;
rom[646] = 32'h6628A0EF;
rom[647] = 32'h090704E3;
rom[648] = 32'h01C7B633;
rom[649] = 32'hDF720B6F;
rom[650] = 32'hAC86A513;
rom[651] = 32'h372D5063;
rom[652] = 32'h00C32103;
rom[653] = 32'hB169A823;
rom[654] = 32'h87A02823;
rom[655] = 32'hCC43AF93;
rom[656] = 32'h01C9AD83;
rom[657] = 32'h010CD893;
rom[658] = 32'h146231EF;
rom[659] = 32'h0103AF83;
rom[660] = 32'h00C0A203;
rom[661] = 32'h01AB3B33;
rom[662] = 32'hF20026EF;
rom[663] = 32'h00FA48B3;
rom[664] = 32'h00C3A183;
rom[665] = 32'h01052503;
rom[666] = 32'h770C0C93;
rom[667] = 32'h012927B3;
rom[668] = 32'h01BDA423;
rom[669] = 32'h000BA603;
rom[670] = 32'hA9CDC86F;
rom[671] = 32'h3F232A23;
rom[672] = 32'h585AA823;
rom[673] = 32'h80CF0F6F;
rom[674] = 32'h59982223;
rom[675] = 32'h35A64BEF;
rom[676] = 32'h859484EF;
rom[677] = 32'h3B888A93;
rom[678] = 32'hCD420A13;
rom[679] = 32'h6E1C9C63;
rom[680] = 32'hF640A223;
rom[681] = 32'h000F2703;
rom[682] = 32'h14806013;
rom[683] = 32'h44802423;
rom[684] = 32'h00C52D83;
rom[685] = 32'h000629B3;
rom[686] = 32'h5829C863;
rom[687] = 32'hCA972A23;
rom[688] = 32'h40489863;
rom[689] = 32'h000A2A83;
rom[690] = 32'hB6AEDD6F;
rom[691] = 32'h00600AB3;
rom[692] = 32'h018AAA03;
rom[693] = 32'h130DC113;
rom[694] = 32'h019C33B3;
rom[695] = 32'h87824693;
rom[696] = 32'h54162E23;
rom[697] = 32'h19F7FC63;
rom[698] = 32'h5F06B4EF;
rom[699] = 32'h178B9C63;
rom[700] = 32'h79817D13;
rom[701] = 32'h4552E463;
rom[702] = 32'h41DED6B3;
rom[703] = 32'h0088A003;
rom[704] = 32'h000F2083;
rom[705] = 32'h428BAE23;
rom[706] = 32'h000BA333;
rom[707] = 32'hA34BE293;
rom[708] = 32'h64B50CE3;
rom[709] = 32'h01E630B3;
rom[710] = 32'hB4602623;
rom[711] = 32'h9D9D7EEF;
rom[712] = 32'h004C7E33;
rom[713] = 32'hF2709E6F;
rom[714] = 32'h002A73B3;
rom[715] = 32'hCD54C76F;
rom[716] = 32'h5E441863;
rom[717] = 32'h000F9BB3;
rom[718] = 32'h408F5C13;
rom[719] = 32'hF5102E23;
rom[720] = 32'h1F011863;
rom[721] = 32'h005FA333;
rom[722] = 32'h012200B3;
rom[723] = 32'h40AF0933;
rom[724] = 32'h4A955C63;
rom[725] = 32'h01C6A283;
rom[726] = 32'h0080A203;
rom[727] = 32'h16AA8463;
rom[728] = 32'h2AFEA623;
rom[729] = 32'h914DAD13;
rom[730] = 32'h011961B3;
rom[731] = 32'hAFF0AA23;
rom[732] = 32'h85CB9013;
rom[733] = 32'hE40B8593;
rom[734] = 32'h6D8DAC13;
rom[735] = 32'h838DF613;
rom[736] = 32'h5902E693;
rom[737] = 32'h2A924A6F;
rom[738] = 32'h6114DCE3;
rom[739] = 32'h01219EB3;
rom[740] = 32'h00D78233;
rom[741] = 32'h411CDFB3;
rom[742] = 32'h2201FD93;
rom[743] = 32'h07672823;
rom[744] = 32'hA9C21193;
rom[745] = 32'h13809D13;
rom[746] = 32'h410A5A13;
rom[747] = 32'h0103A083;
rom[748] = 32'h80A2AA23;
rom[749] = 32'h1F823393;
rom[750] = 32'h01A4B933;
rom[751] = 32'h9FC981EF;
rom[752] = 32'hA1B2A623;
rom[753] = 32'h18859E93;
rom[754] = 32'h11C62223;
rom[755] = 32'hBFE02E23;
rom[756] = 32'h00C42803;
rom[757] = 32'hC6826F13;
rom[758] = 32'h400ADD93;
rom[759] = 32'hAB811993;
rom[760] = 32'h0ED9BDEF;
rom[761] = 32'h051E1063;
rom[762] = 32'hF25CA423;
rom[763] = 32'hF2832823;
rom[764] = 32'h32062C23;
rom[765] = 32'h01C42283;
rom[766] = 32'hA2C4FF13;
rom[767] = 32'h011AC833;
rom[768] = 32'h406E82B3;
rom[769] = 32'hDA9CA223;
rom[770] = 32'h3A248863;
rom[771] = 32'hC7E6AE23;
rom[772] = 32'h01452E83;
rom[773] = 32'h0188DB93;
rom[774] = 32'h9C0B8FEF;
rom[775] = 32'h01462603;
rom[776] = 32'h46823213;
rom[777] = 32'h602DE0EF;
rom[778] = 32'h0045AC83;
rom[779] = 32'hD2C72423;
rom[780] = 32'h6646C593;
rom[781] = 32'h01FD7833;
rom[782] = 32'h501CE063;
rom[783] = 32'hE8E9DC6F;
rom[784] = 32'h0080A683;
rom[785] = 32'h58FB2C23;
rom[786] = 32'h41825E13;
rom[787] = 32'h2B8AA713;
rom[788] = 32'h31171463;
rom[789] = 32'h726A736F;
rom[790] = 32'hAEC60513;
rom[791] = 32'hB02BAE23;
rom[792] = 32'h018EA803;
rom[793] = 32'h01882403;
rom[794] = 32'hAFAF17EF;
rom[795] = 32'h45BFAE23;
rom[796] = 32'h3611D8E3;
rom[797] = 32'h004AD313;
rom[798] = 32'h59D84063;
rom[799] = 32'h0080AD03;
rom[800] = 32'h2F25DF6F;
rom[801] = 32'h01442903;
rom[802] = 32'h1A89A223;
rom[803] = 32'h089B04E3;
rom[804] = 32'h96B4A823;
rom[805] = 32'h4A6480E3;
rom[806] = 32'h0182AA03;
rom[807] = 32'h9BCE4D13;
rom[808] = 32'hE84C4293;
rom[809] = 32'h26F398E3;
rom[810] = 32'hA003BA13;
rom[811] = 32'h1EEA1C63;
rom[812] = 32'h94896B13;
rom[813] = 32'h87CDFF13;
rom[814] = 32'h7AB770E3;
rom[815] = 32'h743860E3;
rom[816] = 32'h69922223;
rom[817] = 32'h4B5B7063;
rom[818] = 32'h25254CEF;
rom[819] = 32'h7049FC13;
rom[820] = 32'hA9252223;
rom[821] = 32'h00042A83;
rom[822] = 32'hE930C76F;
rom[823] = 32'hF360AA23;
rom[824] = 32'h0106A803;
rom[825] = 32'h225C2A23;
rom[826] = 32'h75166A6F;
rom[827] = 32'h76CDF0E3;
rom[828] = 32'h008B2AB3;
rom[829] = 32'hA801B693;
rom[830] = 32'h7B0AA223;
rom[831] = 32'hBB32146F;
rom[832] = 32'h58828993;
rom[833] = 32'hC7C56213;
rom[834] = 32'hA940C393;
rom[835] = 32'hA632A023;
rom[836] = 32'h00C0A983;
rom[837] = 32'h008E2703;
rom[838] = 32'h0F0C1E6F;
rom[839] = 32'h01412703;
rom[840] = 32'hBD078213;
rom[841] = 32'h090CA023;
rom[842] = 32'hC9B9E1EF;
rom[843] = 32'h01F8206F;
rom[844] = 32'h008E2083;
rom[845] = 32'h57729CE3;
rom[846] = 32'h6FEA10E3;
rom[847] = 32'h9CBE2823;
rom[848] = 32'h5B094E13;
rom[849] = 32'h37442423;
rom[850] = 32'h010AAB83;
rom[851] = 32'h628D4863;
rom[852] = 32'h0087AD83;
rom[853] = 32'h004EAA03;
rom[854] = 32'h656014E3;
rom[855] = 32'h1647AE23;
rom[856] = 32'h011DCD33;
rom[857] = 32'h4044DCB3;
rom[858] = 32'h254B1063;
rom[859] = 32'h5CF72623;
rom[860] = 32'h5393ECE3;
rom[861] = 32'hFED7A823;
rom[862] = 32'h3404F8E3;
rom[863] = 32'h330B1613;
rom[864] = 32'h41805D13;
rom[865] = 32'h01042983;
rom[866] = 32'h014AAB03;
rom[867] = 32'h8A182C23;
rom[868] = 32'h41505CB3;
rom[869] = 32'h01C11FB3;
rom[870] = 32'hE685896F;
rom[871] = 32'h00D09233;
rom[872] = 32'h5B032223;
rom[873] = 32'hDCB23AEF;
rom[874] = 32'h0041A203;
rom[875] = 32'h401CA76F;
rom[876] = 32'h000E2F03;
rom[877] = 32'h094A4793;
rom[878] = 32'h9FF4A06F;
rom[879] = 32'h0101D113;
rom[880] = 32'h2E171463;
rom[881] = 32'hC2CD9C13;
rom[882] = 32'h00C04833;
rom[883] = 32'h5DC6F513;
rom[884] = 32'hF67D2E23;
rom[885] = 32'h01542633;
rom[886] = 32'h24682A23;
rom[887] = 32'h0BECD16F;
rom[888] = 32'h33E06D6F;
rom[889] = 32'hE649A623;
rom[890] = 32'h725A9463;
rom[891] = 32'h11912C23;
rom[892] = 32'h06761463;
rom[893] = 32'h296510E3;
rom[894] = 32'h58839E13;
rom[895] = 32'h2E0BAE23;
rom[896] = 32'h01CF2683;
rom[897] = 32'hCE10A623;
rom[898] = 32'h0004A983;
rom[899] = 32'hB9F1486F;
rom[900] = 32'hFB4DA823;
rom[901] = 32'h015CF7B3;
rom[902] = 32'h008E2083;
rom[903] = 32'h97CCF76F;
rom[904] = 32'h8FE59A6F;
rom[905] = 32'h77449113;
rom[906] = 32'h3DCC9E93;
rom[907] = 32'h00C62103;
rom[908] = 32'h198960E3;
rom[909] = 32'h00486133;
rom[910] = 32'hD5F230EF;
rom[911] = 32'hCC8ACF93;
rom[912] = 32'h40CDD693;
rom[913] = 32'h56708463;
rom[914] = 32'h018FD493;
rom[915] = 32'h012A62B3;
rom[916] = 32'h004A2383;
rom[917] = 32'h00AA3F33;
rom[918] = 32'h00B46EB3;
rom[919] = 32'h1F062B6F;
rom[920] = 32'h6ECA266F;
rom[921] = 32'h6803F4E3;
rom[922] = 32'h01CCAB03;
rom[923] = 32'h1D81E193;
rom[924] = 32'hB27A6B6F;
rom[925] = 32'h2FA9CC63;
rom[926] = 32'h7230A023;
rom[927] = 32'h000BA203;
rom[928] = 32'h41CEA823;
rom[929] = 32'h40F65FB3;
rom[930] = 32'h02BB2E23;
rom[931] = 32'h5397EF6F;
rom[932] = 32'h004FAC83;
rom[933] = 32'h015C0433;
rom[934] = 32'h0180AF03;
rom[935] = 32'h01C6A683;
rom[936] = 32'h17EAA823;
rom[937] = 32'h2942BE93;
rom[938] = 32'h0084AD03;
rom[939] = 32'hA32C2823;
rom[940] = 32'h4B56E463;
rom[941] = 32'h5221AE23;
rom[942] = 32'h22C6F8E3;
rom[943] = 32'h9802AA13;
rom[944] = 32'h5F2108E3;
rom[945] = 32'h194790E3;
rom[946] = 32'h0083AF03;
rom[947] = 32'h00C92683;
rom[948] = 32'h325D50EF;
rom[949] = 32'hE56083EF;
rom[950] = 32'h4E0D0863;
rom[951] = 32'h01593BB3;
rom[952] = 32'h0131D9B3;
rom[953] = 32'h15B7F0E3;
rom[954] = 32'h0702FB93;
rom[955] = 32'hB8422223;
rom[956] = 32'h008FB633;
rom[957] = 32'h208F8E93;
rom[958] = 32'h2F97E863;
rom[959] = 32'h4D574CE3;
rom[960] = 32'hF587A423;
rom[961] = 32'hD2B89EEF;
rom[962] = 32'h7A36C063;
rom[963] = 32'hE699266F;
rom[964] = 32'hC79CFD6F;
rom[965] = 32'h29824493;
rom[966] = 32'h9ECF6593;
rom[967] = 32'h2462A823;
rom[968] = 32'h5BE810E3;
rom[969] = 32'h01C4A783;
rom[970] = 32'h0082AE83;
rom[971] = 32'hF5442823;
rom[972] = 32'h70290C63;
rom[973] = 32'hC2CDF713;
rom[974] = 32'h6583E513;
rom[975] = 32'h6F030463;
rom[976] = 32'h01832903;
rom[977] = 32'h28CDCCE3;
rom[978] = 32'h36E8A823;
rom[979] = 32'h0009AC83;
rom[980] = 32'h462BD4E3;
rom[981] = 32'h74F41463;
rom[982] = 32'hDE17A623;
rom[983] = 32'h18EF2223;
rom[984] = 32'h008F5E13;
rom[985] = 32'h22DD9863;
rom[986] = 32'h2CC92423;
rom[987] = 32'h00CC9133;
rom[988] = 32'h0186E433;
rom[989] = 32'hAB8B0D13;
rom[990] = 32'hC4CC1493;
rom[991] = 32'h73A598E3;
rom[992] = 32'h01CE2283;
rom[993] = 32'h8DE0D2EF;
rom[994] = 32'h0089A403;
rom[995] = 32'h110D7C93;
rom[996] = 32'h00CAA503;
rom[997] = 32'h9B1B97EF;
rom[998] = 32'h01CB2803;
rom[999] = 32'h93B82823;
rom[1000] = 32'h5B806463;
rom[1001] = 32'hB1F850EF;
rom[1002] = 32'h4BEFE1EF;
rom[1003] = 32'h5D69D463;
rom[1004] = 32'h01882983;
rom[1005] = 32'h410D5713;
rom[1006] = 32'h41C2D213;
rom[1007] = 32'h00554BB3;
rom[1008] = 32'h43B7F0E3;
rom[1009] = 32'h3F8FC713;
rom[1010] = 32'h2CCC78E3;
rom[1011] = 32'h00CD2E03;
rom[1012] = 32'h7EA940E3;
rom[1013] = 32'h18022E23;
rom[1014] = 32'hE2AF646F;
rom[1015] = 32'hA7012893;
rom[1016] = 32'hEDFE2E23;
rom[1017] = 32'h54328463;
rom[1018] = 32'h7D48D463;
rom[1019] = 32'h39CA94E3;
rom[1020] = 32'h014BE633;
rom[1021] = 32'h0183D893;
rom[1022] = 32'hFF41B093;
rom[1023] = 32'h290114E3;

    end
    // Assign output
    always @(posedge clk) begin
        instr <= rom[addr];
    end
    
endmodule
    